`define BYTE0 0
`define BYTE1 1
`define BYTE2 2
`define BYTE3 3
`define ENABLE 4
`define DISABLE 5
`define SET 6

`define ACK 7
