module sine_lut(addr, s);

input [7:0] addr;
output [7:0] s;

reg [7:0] s;

always @(addr) begin
case (addr)
0: s = 8'h80;
1: s = 8'h83;
2: s = 8'h86;
3: s = 8'h89;
4: s = 8'h8C;
5: s = 8'h8F;
6: s = 8'h92;
7: s = 8'h95;
8: s = 8'h98;
9: s = 8'h9B;
10: s = 8'h9E;
11: s = 8'hA2;
12: s = 8'hA5;
13: s = 8'hA7;
14: s = 8'hAA;
15: s = 8'hAD;
16: s = 8'hB0;
17: s = 8'hB3;
18: s = 8'hB6;
19: s = 8'hB9;
20: s = 8'hBC;
21: s = 8'hBE;
22: s = 8'hC1;
23: s = 8'hC4;
24: s = 8'hC6;
25: s = 8'hC9;
26: s = 8'hCB;
27: s = 8'hCE;
28: s = 8'hD0;
29: s = 8'hD3;
30: s = 8'hD5;
31: s = 8'hD7;
32: s = 8'hDA;
33: s = 8'hDC;
34: s = 8'hDE;
35: s = 8'hE0;
36: s = 8'hE2;
37: s = 8'hE4;
38: s = 8'hE6;
39: s = 8'hE8;
40: s = 8'hEA;
41: s = 8'hEB;
42: s = 8'hED;
43: s = 8'hEE;
44: s = 8'hF0;
45: s = 8'hF1;
46: s = 8'hF3;
47: s = 8'hF4;
48: s = 8'hF5;
49: s = 8'hF6;
50: s = 8'hF8;
51: s = 8'hF9;
52: s = 8'hFA;
53: s = 8'hFA;
54: s = 8'hFB;
55: s = 8'hFC;
56: s = 8'hFD;
57: s = 8'hFD;
58: s = 8'hFE;
59: s = 8'hFE;
60: s = 8'hFE;
61: s = 8'hFF;
62: s = 8'hFF;
63: s = 8'hFF;
64: s = 8'hFF;
65: s = 8'hFF;
66: s = 8'hFF;
67: s = 8'hFF;
68: s = 8'hFE;
69: s = 8'hFE;
70: s = 8'hFE;
71: s = 8'hFD;
72: s = 8'hFD;
73: s = 8'hFC;
74: s = 8'hFB;
75: s = 8'hFA;
76: s = 8'hFA;
77: s = 8'hF9;
78: s = 8'hF8;
79: s = 8'hF6;
80: s = 8'hF5;
81: s = 8'hF4;
82: s = 8'hF3;
83: s = 8'hF1;
84: s = 8'hF0;
85: s = 8'hEE;
86: s = 8'hED;
87: s = 8'hEB;
88: s = 8'hEA;
89: s = 8'hE8;
90: s = 8'hE6;
91: s = 8'hE4;
92: s = 8'hE2;
93: s = 8'hE0;
94: s = 8'hDE;
95: s = 8'hDC;
96: s = 8'hDA;
97: s = 8'hD7;
98: s = 8'hD5;
99: s = 8'hD3;
100: s = 8'hD0;
101: s = 8'hCE;
102: s = 8'hCB;
103: s = 8'hC9;
104: s = 8'hC6;
105: s = 8'hC4;
106: s = 8'hC1;
107: s = 8'hBE;
108: s = 8'hBC;
109: s = 8'hB9;
110: s = 8'hB6;
111: s = 8'hB3;
112: s = 8'hB0;
113: s = 8'hAD;
114: s = 8'hAA;
115: s = 8'hA7;
116: s = 8'hA5;
117: s = 8'hA2;
118: s = 8'h9E;
119: s = 8'h9B;
120: s = 8'h98;
121: s = 8'h95;
122: s = 8'h92;
123: s = 8'h8F;
124: s = 8'h8C;
125: s = 8'h89;
126: s = 8'h86;
127: s = 8'h83;
128: s = 8'h80;
129: s = 8'h7C;
130: s = 8'h79;
131: s = 8'h76;
132: s = 8'h73;
133: s = 8'h70;
134: s = 8'h6D;
135: s = 8'h6A;
136: s = 8'h67;
137: s = 8'h64;
138: s = 8'h61;
139: s = 8'h5D;
140: s = 8'h5A;
141: s = 8'h58;
142: s = 8'h55;
143: s = 8'h52;
144: s = 8'h4F;
145: s = 8'h4C;
146: s = 8'h49;
147: s = 8'h46;
148: s = 8'h43;
149: s = 8'h41;
150: s = 8'h3E;
151: s = 8'h3B;
152: s = 8'h39;
153: s = 8'h36;
154: s = 8'h34;
155: s = 8'h31;
156: s = 8'h2F;
157: s = 8'h2C;
158: s = 8'h2A;
159: s = 8'h28;
160: s = 8'h25;
161: s = 8'h23;
162: s = 8'h21;
163: s = 8'h1F;
164: s = 8'h1D;
165: s = 8'h1B;
166: s = 8'h19;
167: s = 8'h17;
168: s = 8'h15;
169: s = 8'h14;
170: s = 8'h12;
171: s = 8'h11;
172: s = 8'h0F;
173: s = 8'h0E;
174: s = 8'h0C;
175: s = 8'h0B;
176: s = 8'h0A;
177: s = 8'h09;
178: s = 8'h07;
179: s = 8'h06;
180: s = 8'h05;
181: s = 8'h05;
182: s = 8'h04;
183: s = 8'h03;
184: s = 8'h02;
185: s = 8'h02;
186: s = 8'h01;
187: s = 8'h01;
188: s = 8'h01;
189: s = 8'h00;
190: s = 8'h00;
191: s = 8'h00;
192: s = 8'h00;
193: s = 8'h00;
194: s = 8'h00;
195: s = 8'h00;
196: s = 8'h01;
197: s = 8'h01;
198: s = 8'h01;
199: s = 8'h02;
200: s = 8'h02;
201: s = 8'h03;
202: s = 8'h04;
203: s = 8'h05;
204: s = 8'h05;
205: s = 8'h06;
206: s = 8'h07;
207: s = 8'h09;
208: s = 8'h0A;
209: s = 8'h0B;
210: s = 8'h0C;
211: s = 8'h0E;
212: s = 8'h0F;
213: s = 8'h11;
214: s = 8'h12;
215: s = 8'h14;
216: s = 8'h15;
217: s = 8'h17;
218: s = 8'h19;
219: s = 8'h1B;
220: s = 8'h1D;
221: s = 8'h1F;
222: s = 8'h21;
223: s = 8'h23;
224: s = 8'h25;
225: s = 8'h28;
226: s = 8'h2A;
227: s = 8'h2C;
228: s = 8'h2F;
229: s = 8'h31;
230: s = 8'h34;
231: s = 8'h36;
232: s = 8'h39;
233: s = 8'h3B;
234: s = 8'h3E;
235: s = 8'h41;
236: s = 8'h43;
237: s = 8'h46;
238: s = 8'h49;
239: s = 8'h4C;
240: s = 8'h4F;
241: s = 8'h52;
242: s = 8'h55;
243: s = 8'h58;
244: s = 8'h5A;
245: s = 8'h5D;
246: s = 8'h61;
247: s = 8'h64;
248: s = 8'h67;
249: s = 8'h6A;
250: s = 8'h6D;
251: s = 8'h70;
252: s = 8'h73;
253: s = 8'h76;
254: s = 8'h79;
255: s = 8'h7C;
endcase
end
endmodule

